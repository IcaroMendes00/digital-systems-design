// hello world in verilog
module hello_world();
    initial begin
        $display("\n\t Hello World! \n");
    end
endmodule

// task 1
module say_my_name();
    initial begin
        $display("\n\t  My name is Icaro Mendes and I start the course today 4 Jun 2024. \n");
    end
endmodule