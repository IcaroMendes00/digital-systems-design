// manipulacao de vetores em verilog
// exercise 4

module vector_manipulation();

// registradores
    reg [7:0] a = 0; // registrador/vetor de 8bits (MSB = 7, LSB = 0) 
    reg [6:0] b = 0; // registrador/vetor de 7bits 
    reg [7:0] d = 0; // registrador/vetor de 8bits 
// fios
    wire [1:0] c;    // net de 2bits

// procedimentos
// procedimento 1 - atibuicao continua entre o registrador e fio
// c[1] = a[3]
// c[0] = a[2]
    assign c[1:0] = a[3:2]; // 'bit slicing'

// procedimento 2 - verifica continuamente os valores de a, b, c e d
    initial begin
        $monitor("\n\t PROC 2 - a = %b, b = %b, c = %b, d = %b", a, b, c, d);
    end

// procedimento 3 - mudanca de valores
    initial begin
        #1 a = 1;
        #1 a = 8'b1111_0101;
        #1 a = 8'b1111_1000;
        #1 a = 8'b0000_1000;
        #1 a = 8'b0;

        #1 b = 7'b111_1111;
        #1 d[3:0] = a[3:0];
        #1 d[7:4] = b[6:3];

        #1 a = 8'b0000_1110;
        #1 d = {a[3:0], b[3:0]};
        #1 d = {b[3:0], a[7:4]};
    end

endmodule
// end of file